module SYS_CTRL #(parameter WIDTH=8,DEPTH=4) ( input CLK,RST,
                                               input [WIDTH*2-1:0] ALU_OUT,
                                               input OUT_VALID,
                                               input [WIDTH-1:0] RD_DATA,
                                               input RD_DATA_valid,
                                               input [WIDTH-1:0] RX_P_DATA,
                                               input RX_D_VLD,
                                               input FIFO_FULL,
                                               output reg ENABLE,CLK_EN,
                                               output reg [3:0] ALU_FUN,
                                               output reg [DEPTH-1:0] ADDRESS,
                                               output reg WrEn,RdEn,
                                               output reg [WIDTH-1:0] WrData,
                                               output reg [WIDTH-1:0] TX_P_DATA,
                                               output reg TX_D_VLD
                                               );
localparam IDLE=4'b0000,
    DECODE=4'b0001,
    WRITE_ADDR=4'b0010,
    WRITE_DATA=4'b0011,
    READ_ADDR=4'b0100,
    SEND_FIFO=4'b0101,
    ALU_FUNC=4'b0110,
    OPERAND_A=4'b0111,
    OPERAND_B=4'b1000,
    ALU_STORE=4'b1001,
    ALU_FIFO=4'b1010;

reg [3:0] CURRENT_STATE,NEXT_STATE;
reg [DEPTH-1:0] ADDRESS_comp,ADDRESS_reg;
reg ADDR_FLAG,ALU_FLAG;
reg count,count_comp;
reg [2*WIDTH-1:0] ALU_OUT_REG;
always@(posedge CLK, negedge RST)////////current state logic
  begin
    if(!RST)
      begin
        CURRENT_STATE<=IDLE;
        count<=0;
      end
    else
      begin
        CURRENT_STATE<=NEXT_STATE;
        count<=count_comp;
      end
  end

always@(*)
  begin
    NEXT_STATE=IDLE;
    count_comp=0;
    case(CURRENT_STATE)
      IDLE:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=DECODE;
            end
          else
            begin
              NEXT_STATE=IDLE;
            end
        end
      DECODE:
        begin
              case(RX_P_DATA)
                'hAA:
                  begin
                    NEXT_STATE=WRITE_ADDR;
                  end
                'hBB:
                  begin
                    NEXT_STATE=READ_ADDR;
                  end
                'hCC:
                  begin
                    NEXT_STATE=OPERAND_A;
                  end
                'hDD:
                  begin
                    NEXT_STATE=ALU_FUNC;
                  end
                default:
                  begin
                    NEXT_STATE=IDLE;
                  end
              endcase     
        end
      WRITE_ADDR:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=WRITE_DATA;
            end
          else
            begin
              NEXT_STATE=WRITE_ADDR;
            end
        end
      WRITE_DATA:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=IDLE;
            end
          else
            begin
              NEXT_STATE=WRITE_DATA;
            end
        end
      READ_ADDR:
        begin
          if(RD_DATA_valid)
            begin
              NEXT_STATE=SEND_FIFO;
            end
          else
            begin
              NEXT_STATE=READ_ADDR;
            end
        end
      SEND_FIFO:
        begin
          if(FIFO_FULL)
            begin
              NEXT_STATE=SEND_FIFO;
            end
          else
            begin
              if(RX_D_VLD)
                begin
                  NEXT_STATE=DECODE;
                end
              else
                begin
                  NEXT_STATE=IDLE;
                end
            end
        end
      ALU_FUNC:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=ALU_STORE;
            end
          else
            begin
              NEXT_STATE=ALU_FUNC;
            end
        end
      ALU_STORE:
        begin
          if(OUT_VALID)
            begin
              NEXT_STATE=ALU_FIFO;
            end
          else
            begin
              NEXT_STATE=ALU_STORE;
            end
        end
      ALU_FIFO:
        begin
          if(FIFO_FULL)
            begin
              NEXT_STATE=ALU_FIFO;
            end
          else
            if(count)
              begin
                if(RX_D_VLD)
                begin
                  NEXT_STATE=DECODE;
                end
               else
                begin
                  NEXT_STATE=IDLE;
                end
              count_comp=0;
              end
            else
              begin
                NEXT_STATE=ALU_FIFO;
                count_comp=1;
              end
        end
      OPERAND_A:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=OPERAND_B;
            end
          else
            begin
              NEXT_STATE=OPERAND_A;
            end
        end
      OPERAND_B:
        begin
          if(RX_D_VLD)
            begin
              NEXT_STATE=ALU_FUNC;
            end
          else
            begin
              NEXT_STATE=OPERAND_B;
            end
        end
    endcase
  end
  
always@(*)
  begin
    ENABLE=0;
    CLK_EN=0;
    ALU_FUN=0;
    ADDRESS_comp=0;
    ADDR_FLAG=0;
    ADDRESS=0;
    WrEn=0;
    RdEn=0;
    WrData=0;
    TX_P_DATA=0;
    TX_D_VLD=0;
    ALU_FLAG=0;
    case(CURRENT_STATE)
      WRITE_ADDR:
        begin
          if(RX_D_VLD)
            begin
              ADDRESS_comp=RX_P_DATA;
              ADDR_FLAG=1;
            end
          else
            begin
              ADDRESS_comp=0;
              ADDR_FLAG=0;
            end
        end
      WRITE_DATA:
        begin
          if(RX_D_VLD)
            begin
              ADDRESS=ADDRESS_reg;
              WrData=RX_P_DATA;
              WrEn=1;
            end
          else
            begin
              ADDRESS=0;
              WrData=0;
              WrEn=0;
            end
        end
      READ_ADDR:
        begin
          if(RX_D_VLD)
            begin
              RdEn=1;
              ADDRESS=RX_P_DATA;
            end
          else
            begin
             ADDRESS=0;
             RdEn=0; 
            end
        end
      SEND_FIFO:////////////////////
        begin
          if(FIFO_FULL)
            begin
              TX_P_DATA=RD_DATA;
              TX_D_VLD=0;
            end
          else
            begin
              TX_P_DATA=RD_DATA;
              TX_D_VLD=1;
            end
        end
      OPERAND_A:
        begin
          if(RX_D_VLD)
            begin
              ADDRESS='b0;
              WrData=RX_P_DATA;
              WrEn=1;
            end
          else
            begin
              ADDRESS=0;
              WrData=0;
              WrEn=0;
            end
        end
      OPERAND_B:
        begin
          if(RX_D_VLD)
            begin
              ADDRESS='b01;
              WrData=RX_P_DATA;
              WrEn=1;
            end
          else
            begin
              ADDRESS=0;
              WrData=0;
              WrEn=0;
            end
        end
      ALU_FUNC:
        begin
          if(RX_D_VLD)
            begin
              ENABLE=1;
              CLK_EN=1;
              ALU_FUN=RX_P_DATA[3:0];
            end
          else
            begin
              ENABLE=0;
              CLK_EN=0;
              ALU_FUN=RX_P_DATA[3:0];
            end
        end
      ALU_STORE:
        begin
          if(OUT_VALID)
            begin
              ALU_FLAG=1;
            end
          else
            begin
              ALU_FLAG=0;
            end
        end
      ALU_FIFO:
        begin
          if(FIFO_FULL)
            begin
              TX_D_VLD=0;
            end
          else if(count)
            begin
              TX_P_DATA=ALU_OUT_REG[2*WIDTH-1:WIDTH];
              TX_D_VLD=1;
            end
          else
            begin
              TX_P_DATA=ALU_OUT_REG[WIDTH-1:0];
              TX_D_VLD=1;
            end
        end
      default:
        begin
          ENABLE=0;
          CLK_EN=0;
          ALU_FUN=0;
          ADDRESS_comp=0;
          ADDR_FLAG=0;
          WrEn=0;
          RdEn=0;
          WrData=0;
          TX_P_DATA=0;
          TX_D_VLD=0;
          ALU_FLAG=0;
        end
    endcase
  end
always@(posedge CLK,negedge RST)
  begin
    if(!RST)
      begin
        ADDRESS_reg<=0;
      end
    else if(ADDR_FLAG)
      begin
        ADDRESS_reg<=ADDRESS_comp;
      end
  end
  
always@(posedge CLK,negedge RST)
  begin
    if(!RST)
      begin
        ALU_OUT_REG<=0;
      end
    else if(ALU_FLAG)
      begin
        ALU_OUT_REG<=ALU_OUT;
      end
  end  
endmodule

